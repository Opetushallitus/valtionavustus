Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} kl. {{ start-time }} — {{ end-date }} kl. {{ end-time }}

Du kan bearbeta ansökan via denna länk: {{& url }}

Ansökan kan bearbetas ända till  ansökningstidens slut.

Ansökan med redigeringar sparas automatiskt i Utbildningsstyrelsens statsunderstödssystem,
men för att den ska beaktas måste den skickas i väg för behandling innan ansökningstiden tar slut.

OBS! Du kan dela detta meddelande till andra projektpartner, men observera att alla som känner till länken kan bearbeta ansökan.

Mer information om ansökan kan ni få av den ansvariga föredragande (nämns i ansökningsmeddelandet).

Vid tekniska frågor om blanketten kan ni ta kontakt per e-post på adressen statsunderstod@oph.fi.

{{>signature}}
