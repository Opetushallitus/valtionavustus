TODO(sv received)
