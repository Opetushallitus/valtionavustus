[SV] Bästa mottagare,

Ansökan om understöd: {{ avustushaku }}

[SV] Yhteishankkeen {{ register-number }} - {{ project-name }} osapuoli

[SV] Opetushallitus on tarkastanut hankkeen valtionavustusta koskevan loppuselvityksen ja toteaa avustusta koskevan asian käsittelyn päättyneeksi.

[SV] Opetushallitus voi asian käsittelyn päättämisestä huolimatta periä avustuksen tai osan siitä takaisin, jos sen tietoon tulee uusi seikka, joka valtionavustuslain 21 tai 22 §:n mukaisesti velvoittaa tai oikeuttaa takaisinperintään.

{{>signature}}
