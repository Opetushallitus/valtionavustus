Bästa mottagare,

er slutredovisning för användningen av statsunderstödet {{ avustushaku-name }} har ännu inte lämnats in.

Kom ihåg att skicka slutredovisningen för behandling inom utsatt tid, senast {{ loppuselvitys-deadline }}.

Projekt som har beviljats förlängd användningstid för understödet kan ha en sista inlämningsdag för slutredovisningen som avviker från vad som nämns ovan. Den sista inlämningsdagen för redovisningar inom projekt som beviljats förlängd användningstid anges i beslutet som fattats utifrån en ändringsansökan.

Om ett projekt som beviljats förlängd användningstid inte har fått en ny tidsfrist för redovisningen, ska slutredovisningen lämnas in inom två månader efter att den förlängda användningstiden har gått ut.

Länk till er redovisningsblankett: {{& url }}

Mera information får ni vid behov av kontaktpersonen som anges i beslutet. Vid tekniska problem, ta kontakt på adressen valtionavustukset@oph.fi

{{>signature}}
