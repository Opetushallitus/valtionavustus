{{ register-number }} - {{ project-name }}

{{ avustushaku-name }}

Ni kan granska understödsbeslutet via denna länk: {{& url }}

Understödsmottagaren ska följa de villkor och begränsningar som beskrivs i understödsbeslutet och i dess bilagor.

Om ni tar emot understödet i enlighet med beslutet, kan ni påbörja projektet. Understödsbeloppet betalas senast den dag som anges i beslutet.

Om ni inte tar emot understödet i enlighet med beslutet, ska ni meddela om detta till {{^is-jotpa-hakemus}}Utbildningsstyrelsen{{/is-jotpa-hakemus}}{{#is-jotpa-hakemus}}Servicecentret för kontinuerligt lärande och sysselsättning{{/is-jotpa-hakemus}} inom den tidsfrist som anges i beslutet. Anmälan ska göras i statsunderstödssystemet via denna länk: {{& refuse-url }}

{{^include-muutoshaku-link}}Understödsmottagaren ansvarar för att kontaktuppgifterna till den som angetts som kontaktperson i statsunderstödssystemet är uppdaterade. Kontaktpersonen kan bytas ut via länken intill under hela understödets användningstid:{{/include-muutoshaku-link}}
{{#include-muutoshaku-link}}Om det uppstår förändringar som inverkar på användningen av statsunderstödet ska man genast göra en skriftlig ändringsansökan. Man ska framföra tillräckliga motiveringar för ändringarna som ingår i ändringsansökan. I oklara situationer kan understödsmottagaren vara i kontakt med kontaktpersonen som anges i understödsbeslutet innan en ändringsansökan görs.

Understödsmottagaren ansvarar för att kontaktuppgifterna till den person som angetts som kontaktperson i statsunderstödssystemet alltid är uppdaterade. Ni kan göra en ändringsansökan samt byta ut kontaktpersonen och göra ändringar i hens kontaktuppgifter under hela projektperiodens gång via följande länk:{{/include-muutoshaku-link}}
{{& modify-url }}

Begäranden om redovisningar och andra meddelanden som riktas till projektet skickas från adressen {{ from }}. De skickas både till projektets kontaktperson och till den officiella e-postadress som den sökande har angett.

Mottagaren av understöd ska spara detta meddelande och länkarna som ingår i meddelandet.

Vid behov ges närmare information av den person som angetts som kontaktperson i understödsbeslutet.



{{>signature}}
