[SV] Bästa mottagare,

Ansökan om understöd: {{ avustushaku }}

[SV] Yhteishankkeen {{ register-number }} - {{ project-name }} osapuoli

[SV] Olemme vastaanottaneet hankkeen väliselvityksen.

[SV] Väliselvitystä voitte tarkastella tästä linkistä: {{& preview-url }}

[SV] Kun selvitys on käsitelty, ilmoitetaan siitä sähköpostitse avustuksen saajan viralliseen sähköpostiosoitteeseen sekä yhteishankkeen osapuolten yhteyshenkilölle.

{{>signature}}
