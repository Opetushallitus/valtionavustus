Bästa mottagare,

vi har tagit emot er slutredovisning.

{{& hakemus-name }}
{{& register-number }}

Ni kan granska er slutredovisning via denna länk: {{& preview-url }}

Det är möjligt att redigera en redovisning som lämnats in för behandling  via länken i den ursprungliga begäran om redovisning fram till den sista inlämningsdagen för redovisningen. I så fall ska redovisningen inte lämnas in för behandling på nytt, utan ändringarna sparas automatiskt. I logguppgifterna i övre kanten av blanketten kan ni kontrollera att ändringarna har sparats.

Mera information får ni vid behov av kontaktpersonen som anges i ert beslut om understöd. Vid tekniska problem ta kontakt på adressen: valtionavustukset@oph.fi.

Ett e-postmeddelande om att redovisningen har behandlats skickas till understödsmottagarens officiella e-postadress och projektets kontaktperson.
