Bästa mottagare,

ni har en halvfärdig ansökan om statsunderstöd {{ avustushaku-name }}. Observera att ansökningstiden för understödet avslutas {{ paattymispaiva }} kl. {{ paattymisaika }}.

Ansökan och ändringar som görs i ansökan sparas automatiskt i Utbildningsstyrelsens statsunderstödssystem, men för att ansökan ska behandlas behöver den skickas för behandling innan ansökningstiden avslutas. En ansökan som skickats efter att ansökningstiden avslutats kan tas till behandling endast av särskilt vägande skäl.

Ni kommer åt att färdigställa er ansökan via denna länk: {{& url }}

Om ni har beslutat att inte lämna in ansökan föranleder detta meddelande inga åtgärder.