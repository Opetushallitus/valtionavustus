Bästa mottagare,

er ändringsansökan har behandlats.

Projekt: {{ register-number }} - {{ project-name }}

Ni kan granska beslutet via denna länk:
{{& paatos-url }}

Ni kan vid behov göra en ny ändringsansökan via denna länk:
{{& muutoshakemus-url }}

Bilaga: {{ attachment-title }}

Mera information ges vid behov av kontaktpersonen som anges i understödsbeslutet.

Hälsningar,
{{ presenter-name }}

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fornamn.efternamn@oph.fi

