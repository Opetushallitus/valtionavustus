Bästa mottagare,

Ni kan nu fylla i blanketten för slutredovisning för projektet {{ register-number }} "{{ project-name }}".

Blanketten för slutredovisning finns på adressen {{& url }} och den ska lämnas in senast {{ selvitysdate }}.

Med vänlig hälsning

{{ presenter-name }}
Utbildningsstyrelsen

telefon 029 533 1000 (växel)
