Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} klo {{ start-time }} — {{ end-date }} klo {{ end-time }}

Du kan se ansökan via länken: {{& url }}

Mer information ger statsunderstod@oph.fi

Utbildningsstyrelsen
Hagnäskajen 6
PB 380
00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
