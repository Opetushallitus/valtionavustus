Bästa mottagare,

Ni kan nu fylla i blanketten för slutredovisning för projektet {{ register-number }} "{{ project-name }}".

Blanketten för slutredovisning finns på adressen {{& url }} och den ska lämnas in senast {{ selvitysdate }}.

Förutnämnda slutdatum gäller projekt som inte har beviljats förlängning av understödets användningstid. Projekt som har beviljats förlängd användningstid ska bevara den bifogade länken till slutredovisningsblanketten och lämna in slutredovisningen i enlighet med tidtabellen som anges i ändringsbeslutet.

Med vänlig hälsning

{{ presenter-name }}

{{>signature}}
