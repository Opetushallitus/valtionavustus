Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} klo {{ start-time }} — {{ end-date }} klo {{ end-time }}

Du kan se ansökan via länken: {{& url }}

Om du väljer att inte få ett bidrag kan du rapportera det i här länken: {{& refuse-url }}

Anmälan måste skickas senast det datum som anges i beslutet.

Om du ska acceptera det här stöd, måste du gör ingenting.

Den föredragande som ansvarar för ansökningen har nämnts i ansökningsmeddelandet.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380
00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
