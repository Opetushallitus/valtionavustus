Hyvä vastaanottaja,

muutoshakemuksenne on käsitelty.

Hanke: {{ register-number }} - {{ project-name }}

Päätöstä voitte tarkastella tästä linkistä:
{{ & paatos-url }}

Tarvittaessa uuden muutoshakemuksen pääsette tekemään tästä linkistä:
{{ & muutoshakemus-url }}

Liite: {{ attachment-title }

Terveisin,
{{ presenter-name }}

Opetushallitus
Hakaniemenranta 6
PL 380, 00531 Helsinki

puhelin 029 533 1000
etunimi.sukunimi@oph.fi
