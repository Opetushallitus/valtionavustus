Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} kl. {{ start-time }} — {{ end-date }} kl. {{ end-time }}

Du kan bearbeta ansökan via denna länk: {{& url }}

Ansökan kan bearbetas ända till  ansökningstidens slut. Ansökningarna behandlas efter ansökningstiden.

OBS! Du kan dela detta meddelande till andra projektpartner, men observera att de kan också bearbeta ansökan.

Tillägsuppgifter ger statsunderstod@oph.fi

Den föredragande som ansvarar för ansökningen har nämnts i ansökningsmeddelandet.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
