Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} klo {{ start-time }} — {{ end-date }} klo {{ end-time }}

Du kan se ansökan via länken: {{& url }}

Den föredragande som ansvarar för ansökningen har nämnts i ansökningsmeddelandet.

Om du väljer att inte få ett bidrag kan du rapportera det i här länken: {{& refuse-url }}

Utbildningsstyrelsen
Hagnäskajen 6
PB 380
00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
