TODO SV Avustushakemus: {{ avustushaku }}

Hakuaika: {{ start-date }} kl. {{ start-time }} - {{ end-date }} kl. {{ end-time }}

Pääset muokkaamaan avustushakemusta tästä linkistä: {{& url }}

Hakemusta on mahdollista muokata hakuajan loppuun asti. Hakemukset käsitellään hakuajan jälkeen.

Huom! Voit jakaa tämän viestien muille hankkeen kumppaneille, mutta huomaa että
jokainen linkin tietävä voi muokata hakemusta.

Lisätietoja antaa opetusneuvos Leena Koski, puh. 029 533 1106,
sähköposti leena.koski@oph.fi

Opetushallitus
Hakaniemenranta 6
PL 380, 00531 Helsinki

puhelin 029 533 1000
faksi 029 533 1035
etunimi.sukunimi@oph.fi