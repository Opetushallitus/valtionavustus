Statsunderstöd: {{ avustushaku }}

Begäran om komplettering:
"{{ taydennyspyynto }}"

Du kan komplettera ansökan via denna länk: {{& url }}

Ändra endast i de punkter som begäran om komplettering gäller.

Om du har frågor kan vända dig till kontaktpersonen per e-post {{ yhteyshenkilo }}

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors
telefon 029 533 1000
fornamn.efternamn@oph.fi
