Ansökan om understöd: {{ grant-name }}

Er anmälan om att ändra kontaktinformation har lämnats in till Utbildningsstyrelsen.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380
00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
