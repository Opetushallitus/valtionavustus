Ansökning: {{ grant-name }}
Projekt: {{ register-number }} "{{ project-name }}"
Sökande: {{ organization-name }}

Anmälan om ändringen till kontaktuppgifterna har skickats till Utbildningsstyrelsen.

Utbildningsstyrelsen
Hagnäskajen 6,
PB 380, 00531 Helsingfors
