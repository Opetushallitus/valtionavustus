Bästa mottagare,

vi har tagit emot er slutredovisning: {{& preview-url }}

Ni får ett meddelande från adressen no-reply@valtionavustukset.oph.fi, då er slutredovisning har behandlats.

Mera information får ni vid behov av kontaktpersonen som anges i beslutet. Vid tekniska problem, ta kontakt på adressen valtionavustukset@oph.fi
