Bästa mottagare,

er mellanredovisning för användningen av statsunderstödet {{ avustushaku-name }} har ännu inte lämnats in.

Kom ihåg att skicka mellanredovisningen för behandling inom utsatt tid, senast {{ valiselvitys-deadline }}. Länk till er mellanredovisningsblankett: {{& url }}

Mera information får ni vid behov av kontaktpersonen som anges i beslutet. Vid tekniska problem, ta kontakt på adressen valtionavustukset@oph.fi

{{>signature}}
