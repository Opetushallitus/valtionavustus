{{^is-jotpa-hakemus}}
Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors
telefon 029 533 1000
fornamn.efternamn@oph.fi
{{/is-jotpa-hakemus}}
{{#is-jotpa-hakemus}}
Servicecentret för kontinuerligt lärande och sysselsättning
Hagnäskajen 6
PB 380, 00531 Helsingfors
telefon 029 533 1000
fornamn.efternamn@jotpa.fi
{{/is-jotpa-hakemus}}
