Bästa mottagare,

vi har tagit emot er mellanredovisning: {{& valiselvitys-preview-url }}

Ni får ett meddelande från adressen no-reply@valtionavustukset.oph.fi då er mellanredovisning har behandlats.

Mera information får ni vid behov av kontaktpersonen som anges i beslutet. Vid tekniska problem, ta kontakt på adressen valtionavustukset@oph.fi