Ansökan om understöd: {{ grant-name }}

Er anmälan om att ni inte tar emot understödet har lämnats in till {{^is-jotpa-hakemus}}Utbildningsstyrelsen{{/is-jotpa-hakemus}}{{#is-jotpa-hakemus}}Servicecentret för kontinuerligt lärande och sysselsättning{{/is-jotpa-hakemus}}.

{{>signature}}
