Ansökan om understöd: {{ avustushaku }}

Begäran om komplettering:
"{{ change-request }}"

Du kan komplettera ansökan via denna länk: {{& url }}
Ändra bara begärda delar.

Begär tilläggsuppgifter per e-post statsunderstod@oph.fi

Den föredragande som ansvarar för ansökningen har nämnts i ansökningsmeddelandet.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
fornamn.efternamn@ubs.fi
