{{ register-number }} - {{ project-name }}

Ansökan om understöd: {{ avustushaku-name }}

Beslut link: {{& url }}

Om du väljer att inte få ett bidrag kan du rapportera det i här länken: {{& refuse-url }}

Den föredragande som ansvarar för ansökningen har nämnts i beslutet.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fornamn.efternamn@ubs.fi
