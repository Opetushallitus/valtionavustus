[SV] Bästa mottagare,

Ansökan om understöd: {{ avustushaku }}

[SV] Yhteishankkeen {{ register-number }} - {{ project-name }} osapuoli

[SV] Muutoshakemuksenne on käsitelty.

[SV] Päätös muutoshakemukseen: {{& paatos-url }}

[SV] Liitteet: {{ attachment-title }}

[SV] Päähakijayhteisö vastaa yhteydenpidosta Opetushallituksen kanssa.

{{>signature}}
