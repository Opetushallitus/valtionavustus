[SV] Bästa mottagare,

Ansökan om understöd: {{ avustushaku }}

{{ register-number }} - {{ project-name }}

[SV] Päätöstä voitte tarkastella tästä linkistä: {{& url }}

{{>signature}}
