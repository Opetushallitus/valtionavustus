Bästa mottagare

det här meddelandet gäller statsunderstödet: {{& register-number }} {{ project-name }}

Vi har tagit emot kompletteringarna till er slutredovisning och den går nu vidare till nästa skede av granskningen. När slutredovisningen är slutbehandlad sänder vi  ett e-postmeddelande till organisationens officiella e-postadress och kontaktpersonen för mottagaren av statsunderstödet.

Med vänlig hälsning
{{ virkailija-first-name }} {{ virkailija-last-name }}
{{ email-of-virkailija }}