Ansökan om understöd: {{ avustushaku-name }}

Beslut link: {{& url }}

Begär tilläggsuppgifter per e-post statsunderstod@oph.fi

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
fornamn.efternamn@ubs.fi
