[SV] Bästa mottagare,

Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} kl. {{ start-time }} — {{ end-date }} kl. {{ end-time }}

Ni kan granska ansökan via denna länk: {{& url }}

[SV] Hakija voi muokata jo lähetettyä hakemusta alkuperäisen hakemuslinkin kautta hakuajan päättymiseen asti.

[SV] Alkuperäinen hakemuslinkki on toimitettu yhteishankkeen päähakijayhteisön viralliseen sähköpostiosoitteeseen ja yhteyshenkilöille.

[SV] Päähakijayhteisö vastaa yhteydenpidosta Opetushallituksen kanssa.

{{>signature}}
