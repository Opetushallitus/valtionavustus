{{ register-number }} - {{ project-name }}

Ansökan om understöd: {{ avustushaku-name }}

Beslut link: {{& url }}

Den föredragande som ansvarar för ansökningen har nämnts i beslutet.

{{>signature}}
