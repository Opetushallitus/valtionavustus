Bästa mottagare,

Ni kan nu fylla i blanketten för mellanredovisning för projektet {{ register-number }} "{{ project-name }}".

Blanketten för mellanredovisning finns på adressen {{& url }} och den ska lämnas in senast {{ selvitysdate }}.

Med vänlig hälsning

{{ presenter-name }}

{{>signature}}
