{{ register-number }} - {{ project-name }}

Ansökan om understöd: {{ avustushaku-name }}

Beslut link: {{& url }}

Den föredragande som ansvarar för ansökningen har nämnts i beslutet.

{{^is-jotpa-hakemus}}Utbildningsstyrelsen{{/is-jotpa-hakemus}}{{#is-jotpa-hakemus}}Servicecentret för kontinuerligt lärande och sysselsättning{{/is-jotpa-hakemus}}
Hagnäskajen 6
PB 380, 00531 Helsingfors
telefon 029 533 1000
fornamn.efternamn@{{^is-jotpa-hakemus}}oph.fi{{/is-jotpa-hakemus}}{{#is-jotpa-hakemus}}jotpa.fi{{/is-jotpa-hakemus}}
