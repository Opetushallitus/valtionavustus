Ansökning: {{ grant-name }}
Projekt: {{ register-number }} "{{ project-name }}"
Sökande: {{ organization-name }}

Anmälan om ändringen till kontaktuppgifterna har skickats till {{^is-jotpa-hakemus}}Utbildningsstyrelsen{{/is-jotpa-hakemus}}{{#is-jotpa-hakemus}}Servicecentret för kontinuerligt lärande och sysselsättning{{/is-jotpa-hakemus}}.

{{>signature}}
