Bästa mottagare,

vi har tagit emot er slutredovisning.

{{& hakemus-name }}
{{& register-number }}

Ni kan granska er slutredovisning via denna länk: {{& preview-url }}

En slutredovisning som har skickats för behandling kan redigeras via länken till blanketten i den ursprungliga begäran om slutredovisning fram till den sista inlämningsdagen för redovisningen. Om slutredovisningen redigeras ska den inte skickas för behandling på nytt, utan ändringarna sparas automatiskt. I logguppgifterna i övre kanten av blanketten kan ni kontrollera att ändringarna har sparats.

Mera information får ni vid behov av kontaktpersonen som anges i ert beslut om understöd. Vid tekniska problem ta kontakt på adressen: valtionavustukset@oph.fi.

Ett e-postmeddelande om att redovisningen har behandlats skickas till understödsmottagarens officiella e-postadress och projektets kontaktperson.
