Avustushakemus: {{ avustushaku }}

Hakuaika: {{ start-date }} klo {{ start-time }} — {{ end-date }} klo {{ end-time }}

Hakemustanne voitte tarkastella tästä linkistä: {{& url }}

Lisätietoja antaa opetusneuvos Leena Koski, puh. 029 533 1106,
sähköposti leena.koski@oph.fi

Opetushallitus
Hakaniemenranta 6
PL 380, 00531 Helsinki

puhelin 029 533 1000
faksi 029 533 1035
etunimi.sukunimi@oph.fi
