Bästa mottagare,

er ändringsansökan har behandlats.

Projekt: {{ register-number }} - {{ project-name }}

Beslut om ändringsansökan: {{& paatos-url }}

Se tidigare ändringsansökningar och gör vid behov en ny ändringsansökan: {{& muutoshakemus-url }}

Bilaga: {{ attachment-title }}

Mera information ges vid behov av kontaktpersonen som anges i beslutet. 

Hälsningar,
{{ presenter-name }}

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fornamn.efternamn@oph.fi

