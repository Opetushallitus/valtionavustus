{{ register-number }} - {{ project-name }}

Ansökan om understöd: {{ avustushaku-name }}

Beslut link: {{& url }}

Om ni bestämmer er för att inte ta emot understödet kan ni göra en anmälan om detta via denna länk: {{& refuse-url }}

Om ni vill förandra kontaktinformationen kan ni göra en anmälan om detta via denna länk: {{& modify-url }}

Anmälan ska göras senast det datum som framgår ur beslutet.

Om ni tar emot understödet behöver ni inte lämna in någon särskild anmälan om detta.

Den föredragande som ansvarar för ansökningen har nämnts i beslutet.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380, 00531 Helsingfors

telefon 029 533 1000
fornamn.efternamn@ubs.fi
