[SV] Bästa mottagare,

Ansökan om understöd: {{ avustushaku }}

[SV] Yhteishankkeen {{ register-number }} - {{ project-name }} osapuoli

[SV] Avustuspäätöstä voitte tarkastella tästä linkistä: {{& url }}

[SV] Avustuksen saajan tulee noudattaa avustuspäätöksessä sekä sen liitteissä kuvattuja ehtoja ja rajoituksia.

[SV] Yhteishankkeen osapuolten tulee huolehtia siitä, että heidän yhteystietonsa ovat ajan tasalla.

[SV] Yhteishankkeen osapuolten yhteystietojen muutokset päivitetään muutoshakulomakkeella päähakijayhteisön kautta.

[SV] Päähakijayhteisö vastaa yhteydenpidosta Opetushallituksen kanssa.

{{>signature}}
