Ansökan om understöd: {{ avustushaku }}

Ansökningstid: {{ start-date }} klo {{ start-time }} — {{ end-date }} klo {{ end-time }}

Du kan se ansökan via länken: {{& url }}

Den sökande kan via länken uppdatera sin ansökan så länge ansökningstiden pågår. Då ska ansökan ändå inte skickas för behandling på nytt, utan efter att ansökan bearbetats ska man med hjälp av logguppgifterna uppe i hörnet av ansökningsblanketten kontrollera att uppdateringarna har sparats.

Den föredragande som ansvarar för ansökningen har nämnts i ansökningsmeddelandet.

Utbildningsstyrelsen
Hagnäskajen 6
PB 380
00531 Helsingfors

telefon 029 533 1000
fax 029 533 1035
