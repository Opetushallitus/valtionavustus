Hyvä vastaanottaja,

hankkeen {{ register-number }} "{{ project-name }}" väliselvityslomake on nyt täytettävissä.

Väliselvityslomake löytyy osoitteesta {{& url }}, ja se tulee palauttaa {{ valiselvitysdate }} mennessä.

Ystävällisin terveisin

Eevi Esittelijä
Opetushallitus

puhelin 029 533 1000