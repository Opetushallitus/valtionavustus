Hyvä vastaanottaja,

tämä viesti koskee avustusta: {{& register-number }} {{ avustushaku-name }}

Olemme vastaanottaneet loppuselvitystänne koskevat täydennykset ja selvityksenne tarkastus siirtyy seuraavaan vaiheeseen. Kun selvitys on käsitelty, ilmoitetaan siitä sähköpostitse avustuksen saajan viralliseen sähköpostiosoitteeseen sekä yhteyshenkilöille.

Ystävällisin terveisin,
{{ virkailija-first-name }} {{ virkailija-last-name }}
{{ email-of-virkailija }}