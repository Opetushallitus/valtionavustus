Hyvä vastaanottaja,

hankkeen {{ register-number }} "{{ project-name }}" loppuselvityslomake on nyt täytettävissä.

Loppuselvityslomake löytyy osoitteesta {{& url }}, ja se tulee palauttaa {{ selvitysdate }} mennessä.

Ystävällisin terveisin

{{ presenter-name }}
Opetushallitus

puhelin 029 533 1000