Avustushakemus: {{ avustushaku }}

Haku päättyy: {{ end-date }} kl. {{ end-time }}

Pääset muokkaamaan avustushakemusta tästä linkistä: {{& url }}

Huom! Voit jakaa tämän viestien muille hankkeen kumppaneille, mutta huomaa että
jokainen linkin tietävä voi muokata hakemusta.
