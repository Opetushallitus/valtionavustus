Bästa mottagare,

er slutredovisning för användningen av statsunderstödet {{ avustushaku-name }} har ännu inte lämnats in.

Kom ihåg att skicka slutredovisningen för behandling inom utsatt tid, senast {{ loppuselvitysdate }}. Länk till er redovisningsblankett: {{& url }}

Mera information får ni vid behov av kontaktpersonen som anges i beslutet. Vid tekniska problem, ta kontakt på adressen valtionavustukset@oph.fi”.